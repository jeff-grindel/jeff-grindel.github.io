
module adder7_8 ( s, co, a, b, c, d, e, f, g, h, ci );
  output [6:0] s;
  input [6:0] a;
  input [6:0] b;
  input [6:0] c;
  input [6:0] d;
  input [6:0] e;
  input [6:0] f;
  input [6:0] g;
  input [6:0] h;
  input ci;
  output co;
  wire   co1, co2, co3, co4, co5, co6, \a0/c6 , \a0/c5 , \a0/c4 , \a0/c3 ,
         \a0/c2 , \a0/c1 , \a0/a0/n3 , \a0/a0/n2 , \a0/a0/n1 , \a6/c6 ,
         \a6/c5 , \a6/c4 , \a6/c3 , \a6/c2 , \a6/c1 , \a5/c6 , \a5/c5 ,
         \a5/c4 , \a5/c3 , \a5/c2 , \a5/c1 , \a4/c6 , \a4/c5 , \a4/c4 ,
         \a4/c3 , \a4/c2 , \a4/c1 , \a3/c6 , \a3/c5 , \a3/c4 , \a3/c3 ,
         \a3/c2 , \a3/c1 , \a2/c6 , \a2/c5 , \a2/c4 , \a2/c3 , \a2/c2 ,
         \a2/c1 , \a1/c6 , \a1/c5 , \a1/c4 , \a1/c3 , \a1/c2 , \a1/c1 , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193;
  wire   [6:0] s1;
  wire   [6:0] s2;
  wire   [6:0] s3;
  wire   [6:0] s4;
  wire   [6:0] s5;
  wire   [6:0] s6;

  XNOR2X1 \a0/a0/U5  ( .A(a[0]), .B(b[0]), .Y(\a0/a0/n2 ) );
  OAI21X1 \a0/a0/U3  ( .A(\a0/a0/n2 ), .B(\a0/a0/n1 ), .C(n17), .Y(\a0/c1 ) );
  XOR2X1 \a0/a0/U2  ( .A(\a0/a0/n1 ), .B(\a0/a0/n2 ), .Y(s1[0]) );
  XNOR2X1 \a6/a6/U5  ( .A(h[6]), .B(s6[6]), .Y(n192) );
  OAI21X1 \a6/a6/U3  ( .A(n192), .B(n191), .C(n18), .Y(co) );
  XOR2X1 \a6/a6/U2  ( .A(n191), .B(n192), .Y(s[6]) );
  XNOR2X1 \a6/a5/U5  ( .A(h[5]), .B(s6[5]), .Y(n189) );
  OAI21X1 \a6/a5/U3  ( .A(n189), .B(n188), .C(n34), .Y(\a6/c6 ) );
  XOR2X1 \a6/a5/U2  ( .A(n188), .B(n189), .Y(s[5]) );
  XNOR2X1 \a6/a4/U5  ( .A(h[4]), .B(s6[4]), .Y(n186) );
  OAI21X1 \a6/a4/U3  ( .A(n186), .B(n185), .C(n2), .Y(\a6/c5 ) );
  XOR2X1 \a6/a4/U2  ( .A(n185), .B(n186), .Y(s[4]) );
  XNOR2X1 \a6/a3/U5  ( .A(h[3]), .B(s6[3]), .Y(n183) );
  OAI21X1 \a6/a3/U3  ( .A(n183), .B(n182), .C(n19), .Y(\a6/c4 ) );
  XOR2X1 \a6/a3/U2  ( .A(n182), .B(n183), .Y(s[3]) );
  XNOR2X1 \a6/a2/U5  ( .A(h[2]), .B(s6[2]), .Y(n180) );
  OAI21X1 \a6/a2/U3  ( .A(n180), .B(n179), .C(n35), .Y(\a6/c3 ) );
  XOR2X1 \a6/a2/U2  ( .A(n179), .B(n180), .Y(s[2]) );
  XNOR2X1 \a6/a1/U5  ( .A(h[1]), .B(s6[1]), .Y(n177) );
  OAI21X1 \a6/a1/U3  ( .A(n177), .B(n176), .C(n3), .Y(\a6/c2 ) );
  XOR2X1 \a6/a1/U2  ( .A(n176), .B(n177), .Y(s[1]) );
  XNOR2X1 \a6/a0/U5  ( .A(h[0]), .B(s6[0]), .Y(n174) );
  OAI21X1 \a6/a0/U3  ( .A(n174), .B(n173), .C(n20), .Y(\a6/c1 ) );
  XOR2X1 \a6/a0/U2  ( .A(n173), .B(n174), .Y(s[0]) );
  XNOR2X1 \a5/a6/U5  ( .A(g[6]), .B(s5[6]), .Y(n171) );
  OAI21X1 \a5/a6/U3  ( .A(n171), .B(n170), .C(n36), .Y(co6) );
  XOR2X1 \a5/a6/U2  ( .A(n170), .B(n171), .Y(s6[6]) );
  XNOR2X1 \a5/a5/U5  ( .A(g[5]), .B(s5[5]), .Y(n168) );
  OAI21X1 \a5/a5/U3  ( .A(n168), .B(n167), .C(n4), .Y(\a5/c6 ) );
  XOR2X1 \a5/a5/U2  ( .A(n167), .B(n168), .Y(s6[5]) );
  XNOR2X1 \a5/a4/U5  ( .A(g[4]), .B(s5[4]), .Y(n165) );
  OAI21X1 \a5/a4/U3  ( .A(n165), .B(n164), .C(n21), .Y(\a5/c5 ) );
  XOR2X1 \a5/a4/U2  ( .A(n164), .B(n165), .Y(s6[4]) );
  XNOR2X1 \a5/a3/U5  ( .A(g[3]), .B(s5[3]), .Y(n162) );
  OAI21X1 \a5/a3/U3  ( .A(n162), .B(n161), .C(n37), .Y(\a5/c4 ) );
  XOR2X1 \a5/a3/U2  ( .A(n161), .B(n162), .Y(s6[3]) );
  XNOR2X1 \a5/a2/U5  ( .A(g[2]), .B(s5[2]), .Y(n159) );
  OAI21X1 \a5/a2/U3  ( .A(n159), .B(n158), .C(n5), .Y(\a5/c3 ) );
  XOR2X1 \a5/a2/U2  ( .A(n158), .B(n159), .Y(s6[2]) );
  XNOR2X1 \a5/a1/U5  ( .A(g[1]), .B(s5[1]), .Y(n156) );
  OAI21X1 \a5/a1/U3  ( .A(n156), .B(n155), .C(n22), .Y(\a5/c2 ) );
  XOR2X1 \a5/a1/U2  ( .A(n155), .B(n156), .Y(s6[1]) );
  XNOR2X1 \a5/a0/U5  ( .A(g[0]), .B(s5[0]), .Y(n153) );
  OAI21X1 \a5/a0/U3  ( .A(n153), .B(n152), .C(n38), .Y(\a5/c1 ) );
  XOR2X1 \a5/a0/U2  ( .A(n152), .B(n153), .Y(s6[0]) );
  XNOR2X1 \a4/a6/U5  ( .A(f[6]), .B(s4[6]), .Y(n150) );
  OAI21X1 \a4/a6/U3  ( .A(n150), .B(n149), .C(n6), .Y(co5) );
  XOR2X1 \a4/a6/U2  ( .A(n149), .B(n150), .Y(s5[6]) );
  XNOR2X1 \a4/a5/U5  ( .A(f[5]), .B(s4[5]), .Y(n147) );
  OAI21X1 \a4/a5/U3  ( .A(n147), .B(n146), .C(n23), .Y(\a4/c6 ) );
  XOR2X1 \a4/a5/U2  ( .A(n146), .B(n147), .Y(s5[5]) );
  XNOR2X1 \a4/a4/U5  ( .A(f[4]), .B(s4[4]), .Y(n144) );
  OAI21X1 \a4/a4/U3  ( .A(n144), .B(n143), .C(n39), .Y(\a4/c5 ) );
  XOR2X1 \a4/a4/U2  ( .A(n143), .B(n144), .Y(s5[4]) );
  XNOR2X1 \a4/a3/U5  ( .A(f[3]), .B(s4[3]), .Y(n141) );
  OAI21X1 \a4/a3/U3  ( .A(n141), .B(n140), .C(n7), .Y(\a4/c4 ) );
  XOR2X1 \a4/a3/U2  ( .A(n140), .B(n141), .Y(s5[3]) );
  XNOR2X1 \a4/a2/U5  ( .A(f[2]), .B(s4[2]), .Y(n138) );
  OAI21X1 \a4/a2/U3  ( .A(n138), .B(n137), .C(n24), .Y(\a4/c3 ) );
  XOR2X1 \a4/a2/U2  ( .A(n137), .B(n138), .Y(s5[2]) );
  XNOR2X1 \a4/a1/U5  ( .A(f[1]), .B(s4[1]), .Y(n135) );
  OAI21X1 \a4/a1/U3  ( .A(n135), .B(n134), .C(n40), .Y(\a4/c2 ) );
  XOR2X1 \a4/a1/U2  ( .A(n134), .B(n135), .Y(s5[1]) );
  XNOR2X1 \a4/a0/U5  ( .A(f[0]), .B(s4[0]), .Y(n132) );
  OAI21X1 \a4/a0/U3  ( .A(n132), .B(n131), .C(n8), .Y(\a4/c1 ) );
  XOR2X1 \a4/a0/U2  ( .A(n131), .B(n132), .Y(s5[0]) );
  XNOR2X1 \a3/a6/U5  ( .A(e[6]), .B(s3[6]), .Y(n129) );
  OAI21X1 \a3/a6/U3  ( .A(n129), .B(n128), .C(n25), .Y(co4) );
  XOR2X1 \a3/a6/U2  ( .A(n128), .B(n129), .Y(s4[6]) );
  XNOR2X1 \a3/a5/U5  ( .A(e[5]), .B(s3[5]), .Y(n126) );
  OAI21X1 \a3/a5/U3  ( .A(n126), .B(n125), .C(n41), .Y(\a3/c6 ) );
  XOR2X1 \a3/a5/U2  ( .A(n125), .B(n126), .Y(s4[5]) );
  XNOR2X1 \a3/a4/U5  ( .A(e[4]), .B(s3[4]), .Y(n123) );
  OAI21X1 \a3/a4/U3  ( .A(n123), .B(n122), .C(n9), .Y(\a3/c5 ) );
  XOR2X1 \a3/a4/U2  ( .A(n122), .B(n123), .Y(s4[4]) );
  XNOR2X1 \a3/a3/U5  ( .A(e[3]), .B(s3[3]), .Y(n120) );
  OAI21X1 \a3/a3/U3  ( .A(n120), .B(n119), .C(n26), .Y(\a3/c4 ) );
  XOR2X1 \a3/a3/U2  ( .A(n119), .B(n120), .Y(s4[3]) );
  XNOR2X1 \a3/a2/U5  ( .A(e[2]), .B(s3[2]), .Y(n117) );
  OAI21X1 \a3/a2/U3  ( .A(n117), .B(n116), .C(n42), .Y(\a3/c3 ) );
  XOR2X1 \a3/a2/U2  ( .A(n116), .B(n117), .Y(s4[2]) );
  XNOR2X1 \a3/a1/U5  ( .A(e[1]), .B(s3[1]), .Y(n114) );
  OAI21X1 \a3/a1/U3  ( .A(n114), .B(n113), .C(n10), .Y(\a3/c2 ) );
  XOR2X1 \a3/a1/U2  ( .A(n113), .B(n114), .Y(s4[1]) );
  XNOR2X1 \a3/a0/U5  ( .A(e[0]), .B(s3[0]), .Y(n111) );
  OAI21X1 \a3/a0/U3  ( .A(n111), .B(n110), .C(n27), .Y(\a3/c1 ) );
  XOR2X1 \a3/a0/U2  ( .A(n110), .B(n111), .Y(s4[0]) );
  XNOR2X1 \a2/a6/U5  ( .A(d[6]), .B(s2[6]), .Y(n108) );
  OAI21X1 \a2/a6/U3  ( .A(n108), .B(n107), .C(n43), .Y(co3) );
  XOR2X1 \a2/a6/U2  ( .A(n107), .B(n108), .Y(s3[6]) );
  XNOR2X1 \a2/a5/U5  ( .A(d[5]), .B(s2[5]), .Y(n105) );
  OAI21X1 \a2/a5/U3  ( .A(n105), .B(n104), .C(n11), .Y(\a2/c6 ) );
  XOR2X1 \a2/a5/U2  ( .A(n104), .B(n105), .Y(s3[5]) );
  XNOR2X1 \a2/a4/U5  ( .A(d[4]), .B(s2[4]), .Y(n102) );
  OAI21X1 \a2/a4/U3  ( .A(n102), .B(n101), .C(n28), .Y(\a2/c5 ) );
  XOR2X1 \a2/a4/U2  ( .A(n101), .B(n102), .Y(s3[4]) );
  XNOR2X1 \a2/a3/U5  ( .A(d[3]), .B(s2[3]), .Y(n99) );
  OAI21X1 \a2/a3/U3  ( .A(n99), .B(n98), .C(n44), .Y(\a2/c4 ) );
  XOR2X1 \a2/a3/U2  ( .A(n98), .B(n99), .Y(s3[3]) );
  XNOR2X1 \a2/a2/U5  ( .A(d[2]), .B(s2[2]), .Y(n96) );
  OAI21X1 \a2/a2/U3  ( .A(n96), .B(n95), .C(n12), .Y(\a2/c3 ) );
  XOR2X1 \a2/a2/U2  ( .A(n95), .B(n96), .Y(s3[2]) );
  XNOR2X1 \a2/a1/U5  ( .A(d[1]), .B(s2[1]), .Y(n93) );
  OAI21X1 \a2/a1/U3  ( .A(n93), .B(n92), .C(n29), .Y(\a2/c2 ) );
  XOR2X1 \a2/a1/U2  ( .A(n92), .B(n93), .Y(s3[1]) );
  XNOR2X1 \a2/a0/U5  ( .A(d[0]), .B(s2[0]), .Y(n90) );
  OAI21X1 \a2/a0/U3  ( .A(n90), .B(n89), .C(n45), .Y(\a2/c1 ) );
  XOR2X1 \a2/a0/U2  ( .A(n89), .B(n90), .Y(s3[0]) );
  XNOR2X1 \a1/a6/U5  ( .A(c[6]), .B(s1[6]), .Y(n87) );
  OAI21X1 \a1/a6/U3  ( .A(n87), .B(n86), .C(n13), .Y(co2) );
  XOR2X1 \a1/a6/U2  ( .A(n86), .B(n87), .Y(s2[6]) );
  XNOR2X1 \a1/a5/U5  ( .A(c[5]), .B(s1[5]), .Y(n84) );
  OAI21X1 \a1/a5/U3  ( .A(n84), .B(n83), .C(n30), .Y(\a1/c6 ) );
  XOR2X1 \a1/a5/U2  ( .A(n83), .B(n84), .Y(s2[5]) );
  XNOR2X1 \a1/a4/U5  ( .A(c[4]), .B(s1[4]), .Y(n81) );
  OAI21X1 \a1/a4/U3  ( .A(n81), .B(n80), .C(n46), .Y(\a1/c5 ) );
  XOR2X1 \a1/a4/U2  ( .A(n80), .B(n81), .Y(s2[4]) );
  XNOR2X1 \a1/a3/U5  ( .A(c[3]), .B(s1[3]), .Y(n78) );
  OAI21X1 \a1/a3/U3  ( .A(n78), .B(n77), .C(n14), .Y(\a1/c4 ) );
  XOR2X1 \a1/a3/U2  ( .A(n77), .B(n78), .Y(s2[3]) );
  XNOR2X1 \a1/a2/U5  ( .A(c[2]), .B(s1[2]), .Y(n75) );
  OAI21X1 \a1/a2/U3  ( .A(n75), .B(n74), .C(n31), .Y(\a1/c3 ) );
  XOR2X1 \a1/a2/U2  ( .A(n74), .B(n75), .Y(s2[2]) );
  XNOR2X1 \a1/a1/U5  ( .A(c[1]), .B(s1[1]), .Y(n72) );
  OAI21X1 \a1/a1/U3  ( .A(n72), .B(n71), .C(n47), .Y(\a1/c2 ) );
  XOR2X1 \a1/a1/U2  ( .A(n71), .B(n72), .Y(s2[1]) );
  XNOR2X1 \a1/a0/U5  ( .A(c[0]), .B(s1[0]), .Y(n69) );
  OAI21X1 \a1/a0/U3  ( .A(n69), .B(n68), .C(n15), .Y(\a1/c1 ) );
  XOR2X1 \a1/a0/U2  ( .A(n68), .B(n69), .Y(s2[0]) );
  XNOR2X1 \a0/a6/U5  ( .A(a[6]), .B(b[6]), .Y(n66) );
  OAI21X1 \a0/a6/U3  ( .A(n66), .B(n65), .C(n32), .Y(co1) );
  XOR2X1 \a0/a6/U2  ( .A(n65), .B(n66), .Y(s1[6]) );
  XNOR2X1 \a0/a5/U5  ( .A(a[5]), .B(b[5]), .Y(n63) );
  OAI21X1 \a0/a5/U3  ( .A(n63), .B(n62), .C(n48), .Y(\a0/c6 ) );
  XOR2X1 \a0/a5/U2  ( .A(n62), .B(n63), .Y(s1[5]) );
  XNOR2X1 \a0/a4/U5  ( .A(a[4]), .B(b[4]), .Y(n60) );
  OAI21X1 \a0/a4/U3  ( .A(n60), .B(n59), .C(n16), .Y(\a0/c5 ) );
  XOR2X1 \a0/a4/U2  ( .A(n59), .B(n60), .Y(s1[4]) );
  XNOR2X1 \a0/a3/U5  ( .A(a[3]), .B(b[3]), .Y(n57) );
  OAI21X1 \a0/a3/U3  ( .A(n57), .B(n56), .C(n33), .Y(\a0/c4 ) );
  XOR2X1 \a0/a3/U2  ( .A(n56), .B(n57), .Y(s1[3]) );
  XNOR2X1 \a0/a2/U5  ( .A(a[2]), .B(b[2]), .Y(n54) );
  OAI21X1 \a0/a2/U3  ( .A(n54), .B(n53), .C(n49), .Y(\a0/c3 ) );
  XOR2X1 \a0/a2/U2  ( .A(n53), .B(n54), .Y(s1[2]) );
  XNOR2X1 \a0/a1/U5  ( .A(a[1]), .B(b[1]), .Y(n51) );
  OAI21X1 \a0/a1/U3  ( .A(n51), .B(n50), .C(n1), .Y(\a0/c2 ) );
  XOR2X1 \a0/a1/U2  ( .A(n50), .B(n51), .Y(s1[1]) );
  AND2X1 U1 ( .A(a[1]), .B(b[1]), .Y(n52) );
  INVX1 U2 ( .A(n52), .Y(n1) );
  AND2X1 U3 ( .A(h[4]), .B(s6[4]), .Y(n187) );
  INVX1 U4 ( .A(n187), .Y(n2) );
  AND2X1 U5 ( .A(h[1]), .B(s6[1]), .Y(n178) );
  INVX1 U6 ( .A(n178), .Y(n3) );
  AND2X1 U7 ( .A(g[5]), .B(s5[5]), .Y(n169) );
  INVX1 U8 ( .A(n169), .Y(n4) );
  AND2X1 U9 ( .A(g[2]), .B(s5[2]), .Y(n160) );
  INVX1 U10 ( .A(n160), .Y(n5) );
  AND2X1 U11 ( .A(f[6]), .B(s4[6]), .Y(n151) );
  INVX1 U12 ( .A(n151), .Y(n6) );
  AND2X1 U13 ( .A(f[3]), .B(s4[3]), .Y(n142) );
  INVX1 U14 ( .A(n142), .Y(n7) );
  AND2X1 U15 ( .A(f[0]), .B(s4[0]), .Y(n133) );
  INVX1 U16 ( .A(n133), .Y(n8) );
  AND2X1 U17 ( .A(e[4]), .B(s3[4]), .Y(n124) );
  INVX1 U18 ( .A(n124), .Y(n9) );
  AND2X1 U19 ( .A(e[1]), .B(s3[1]), .Y(n115) );
  INVX1 U20 ( .A(n115), .Y(n10) );
  AND2X1 U21 ( .A(d[5]), .B(s2[5]), .Y(n106) );
  INVX1 U22 ( .A(n106), .Y(n11) );
  AND2X1 U23 ( .A(d[2]), .B(s2[2]), .Y(n97) );
  INVX1 U24 ( .A(n97), .Y(n12) );
  AND2X1 U25 ( .A(c[6]), .B(s1[6]), .Y(n88) );
  INVX1 U26 ( .A(n88), .Y(n13) );
  AND2X1 U27 ( .A(c[3]), .B(s1[3]), .Y(n79) );
  INVX1 U28 ( .A(n79), .Y(n14) );
  AND2X1 U29 ( .A(c[0]), .B(s1[0]), .Y(n70) );
  INVX1 U30 ( .A(n70), .Y(n15) );
  AND2X1 U31 ( .A(a[4]), .B(b[4]), .Y(n61) );
  INVX1 U32 ( .A(n61), .Y(n16) );
  AND2X1 U33 ( .A(a[0]), .B(b[0]), .Y(\a0/a0/n3 ) );
  INVX1 U34 ( .A(\a0/a0/n3 ), .Y(n17) );
  AND2X1 U35 ( .A(h[6]), .B(s6[6]), .Y(n193) );
  INVX1 U36 ( .A(n193), .Y(n18) );
  AND2X1 U37 ( .A(h[3]), .B(s6[3]), .Y(n184) );
  INVX1 U38 ( .A(n184), .Y(n19) );
  AND2X1 U39 ( .A(h[0]), .B(s6[0]), .Y(n175) );
  INVX1 U40 ( .A(n175), .Y(n20) );
  AND2X1 U41 ( .A(g[4]), .B(s5[4]), .Y(n166) );
  INVX1 U42 ( .A(n166), .Y(n21) );
  AND2X1 U43 ( .A(g[1]), .B(s5[1]), .Y(n157) );
  INVX1 U44 ( .A(n157), .Y(n22) );
  AND2X1 U45 ( .A(f[5]), .B(s4[5]), .Y(n148) );
  INVX1 U46 ( .A(n148), .Y(n23) );
  AND2X1 U47 ( .A(f[2]), .B(s4[2]), .Y(n139) );
  INVX1 U48 ( .A(n139), .Y(n24) );
  AND2X1 U49 ( .A(e[6]), .B(s3[6]), .Y(n130) );
  INVX1 U50 ( .A(n130), .Y(n25) );
  AND2X1 U51 ( .A(e[3]), .B(s3[3]), .Y(n121) );
  INVX1 U52 ( .A(n121), .Y(n26) );
  AND2X1 U53 ( .A(e[0]), .B(s3[0]), .Y(n112) );
  INVX1 U54 ( .A(n112), .Y(n27) );
  AND2X1 U55 ( .A(d[4]), .B(s2[4]), .Y(n103) );
  INVX1 U56 ( .A(n103), .Y(n28) );
  AND2X1 U57 ( .A(d[1]), .B(s2[1]), .Y(n94) );
  INVX1 U58 ( .A(n94), .Y(n29) );
  AND2X1 U59 ( .A(c[5]), .B(s1[5]), .Y(n85) );
  INVX1 U60 ( .A(n85), .Y(n30) );
  AND2X1 U61 ( .A(c[2]), .B(s1[2]), .Y(n76) );
  INVX1 U62 ( .A(n76), .Y(n31) );
  AND2X1 U63 ( .A(a[6]), .B(b[6]), .Y(n67) );
  INVX1 U64 ( .A(n67), .Y(n32) );
  AND2X1 U65 ( .A(a[3]), .B(b[3]), .Y(n58) );
  INVX1 U66 ( .A(n58), .Y(n33) );
  AND2X1 U67 ( .A(h[5]), .B(s6[5]), .Y(n190) );
  INVX1 U68 ( .A(n190), .Y(n34) );
  AND2X1 U69 ( .A(h[2]), .B(s6[2]), .Y(n181) );
  INVX1 U70 ( .A(n181), .Y(n35) );
  AND2X1 U71 ( .A(g[6]), .B(s5[6]), .Y(n172) );
  INVX1 U72 ( .A(n172), .Y(n36) );
  AND2X1 U73 ( .A(g[3]), .B(s5[3]), .Y(n163) );
  INVX1 U74 ( .A(n163), .Y(n37) );
  AND2X1 U75 ( .A(g[0]), .B(s5[0]), .Y(n154) );
  INVX1 U76 ( .A(n154), .Y(n38) );
  AND2X1 U77 ( .A(f[4]), .B(s4[4]), .Y(n145) );
  INVX1 U78 ( .A(n145), .Y(n39) );
  AND2X1 U79 ( .A(f[1]), .B(s4[1]), .Y(n136) );
  INVX1 U80 ( .A(n136), .Y(n40) );
  AND2X1 U81 ( .A(e[5]), .B(s3[5]), .Y(n127) );
  INVX1 U82 ( .A(n127), .Y(n41) );
  AND2X1 U83 ( .A(e[2]), .B(s3[2]), .Y(n118) );
  INVX1 U84 ( .A(n118), .Y(n42) );
  AND2X1 U85 ( .A(d[6]), .B(s2[6]), .Y(n109) );
  INVX1 U86 ( .A(n109), .Y(n43) );
  AND2X1 U87 ( .A(d[3]), .B(s2[3]), .Y(n100) );
  INVX1 U88 ( .A(n100), .Y(n44) );
  AND2X1 U89 ( .A(d[0]), .B(s2[0]), .Y(n91) );
  INVX1 U90 ( .A(n91), .Y(n45) );
  AND2X1 U91 ( .A(c[4]), .B(s1[4]), .Y(n82) );
  INVX1 U92 ( .A(n82), .Y(n46) );
  AND2X1 U93 ( .A(c[1]), .B(s1[1]), .Y(n73) );
  INVX1 U94 ( .A(n73), .Y(n47) );
  AND2X1 U95 ( .A(a[5]), .B(b[5]), .Y(n64) );
  INVX1 U96 ( .A(n64), .Y(n48) );
  AND2X1 U97 ( .A(a[2]), .B(b[2]), .Y(n55) );
  INVX1 U98 ( .A(n55), .Y(n49) );
  INVX2 U99 ( .A(\a0/c2 ), .Y(n53) );
  INVX1 U100 ( .A(\a3/c1 ), .Y(n113) );
  INVX1 U101 ( .A(\a3/c2 ), .Y(n116) );
  INVX1 U102 ( .A(\a3/c3 ), .Y(n119) );
  INVX1 U103 ( .A(\a3/c4 ), .Y(n122) );
  INVX1 U104 ( .A(\a3/c5 ), .Y(n125) );
  INVX1 U105 ( .A(\a0/c1 ), .Y(n50) );
  INVX1 U106 ( .A(\a0/c3 ), .Y(n56) );
  INVX1 U107 ( .A(\a0/c4 ), .Y(n59) );
  INVX1 U108 ( .A(\a0/c5 ), .Y(n62) );
  INVX1 U109 ( .A(\a0/c6 ), .Y(n65) );
  INVX1 U110 ( .A(co1), .Y(n68) );
  INVX1 U111 ( .A(\a1/c1 ), .Y(n71) );
  INVX1 U112 ( .A(\a1/c2 ), .Y(n74) );
  INVX1 U113 ( .A(\a1/c3 ), .Y(n77) );
  INVX1 U114 ( .A(\a1/c4 ), .Y(n80) );
  INVX1 U115 ( .A(\a1/c5 ), .Y(n83) );
  INVX1 U116 ( .A(\a1/c6 ), .Y(n86) );
  INVX1 U117 ( .A(co2), .Y(n89) );
  INVX1 U118 ( .A(\a2/c1 ), .Y(n92) );
  INVX1 U119 ( .A(\a2/c2 ), .Y(n95) );
  INVX1 U120 ( .A(\a2/c3 ), .Y(n98) );
  INVX1 U121 ( .A(\a2/c4 ), .Y(n101) );
  INVX1 U122 ( .A(\a2/c5 ), .Y(n104) );
  INVX1 U123 ( .A(\a2/c6 ), .Y(n107) );
  INVX1 U124 ( .A(co3), .Y(n110) );
  INVX1 U125 ( .A(\a3/c6 ), .Y(n128) );
  INVX1 U126 ( .A(co4), .Y(n131) );
  INVX1 U127 ( .A(\a4/c1 ), .Y(n134) );
  INVX1 U128 ( .A(\a4/c2 ), .Y(n137) );
  INVX1 U129 ( .A(\a4/c3 ), .Y(n140) );
  INVX1 U130 ( .A(\a4/c4 ), .Y(n143) );
  INVX1 U131 ( .A(\a4/c5 ), .Y(n146) );
  INVX1 U132 ( .A(\a4/c6 ), .Y(n149) );
  INVX1 U133 ( .A(co5), .Y(n152) );
  INVX1 U134 ( .A(\a5/c1 ), .Y(n155) );
  INVX1 U135 ( .A(\a5/c2 ), .Y(n158) );
  INVX1 U136 ( .A(\a5/c3 ), .Y(n161) );
  INVX1 U137 ( .A(\a5/c4 ), .Y(n164) );
  INVX1 U138 ( .A(\a5/c5 ), .Y(n167) );
  INVX1 U139 ( .A(\a5/c6 ), .Y(n170) );
  INVX1 U140 ( .A(co6), .Y(n173) );
  INVX1 U141 ( .A(\a6/c1 ), .Y(n176) );
  INVX1 U142 ( .A(\a6/c2 ), .Y(n179) );
  INVX1 U143 ( .A(\a6/c3 ), .Y(n182) );
  INVX1 U144 ( .A(\a6/c4 ), .Y(n185) );
  INVX1 U145 ( .A(\a6/c5 ), .Y(n188) );
  INVX1 U146 ( .A(\a6/c6 ), .Y(n191) );
  INVX1 U147 ( .A(ci), .Y(\a0/a0/n1 ) );
endmodule

