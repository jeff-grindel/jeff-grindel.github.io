
module adder_tree ( s, co, a, b, c, d, e, f, g, h, ci );
  output [6:0] s;
  input [6:0] a;
  input [6:0] b;
  input [6:0] c;
  input [6:0] d;
  input [6:0] e;
  input [6:0] f;
  input [6:0] g;
  input [6:0] h;
  input ci;
  output co;
  wire   \ts2[6] , \a1/ts[6] , \a1/ts[5] , \a1/ts[4] , \a1/ts[3] , \a1/ts[2] ,
         \a1/ts[1] , \a1/ts[0] , \a1/tc[6] , \a1/tc[5] , \a1/tc[4] ,
         \a1/tc[3] , \a1/tc[2] , \a1/tc[1] , \a4/c6 , \a4/c5 , \a4/c4 ,
         \a4/c3 , \a1/s00/n3 , \a1/s00/n2 , \a1/s00/n1 , \a3/ts[6] ,
         \a3/ts[5] , \a3/ts[4] , \a3/ts[3] , \a3/ts[2] , \a3/ts[1] ,
         \a3/tc[6] , \a3/tc[5] , \a3/tc[4] , \a3/tc[3] , \a3/tc[2] ,
         \a2/ts[6] , \a2/ts[5] , \a2/ts[4] , \a2/ts[3] , \a2/ts[2] ,
         \a2/ts[1] , \a2/ts[0] , \a2/tc[6] , \a2/tc[5] , \a2/tc[4] ,
         \a2/tc[3] , \a2/tc[2] , \a2/tc[1] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160;
  wire   [6:0] ts1;
  wire   [6:0] tc1;
  wire   [6:0] tc2;
  wire   [6:0] ts3;
  wire   [6:0] tc3;

  XNOR2X1 \a1/s00/U5  ( .A(a[0]), .B(b[0]), .Y(\a1/s00/n2 ) );
  OAI21X1 \a1/s00/U3  ( .A(\a1/s00/n2 ), .B(\a1/s00/n1 ), .C(n39), .Y(
        \a1/tc[1] ) );
  XOR2X1 \a1/s00/U2  ( .A(\a1/s00/n1 ), .B(\a1/s00/n2 ), .Y(\a1/ts[0] ) );
  XNOR2X1 \a4/a6/U5  ( .A(ts3[6]), .B(tc3[6]), .Y(n159) );
  OAI21X1 \a4/a6/U3  ( .A(n159), .B(n158), .C(n5), .Y(co) );
  XOR2X1 \a4/a6/U2  ( .A(n158), .B(n159), .Y(s[6]) );
  XNOR2X1 \a4/a5/U5  ( .A(ts3[5]), .B(tc3[5]), .Y(n156) );
  OAI21X1 \a4/a5/U3  ( .A(n156), .B(n155), .C(n4), .Y(\a4/c6 ) );
  XOR2X1 \a4/a5/U2  ( .A(n155), .B(n156), .Y(s[5]) );
  XNOR2X1 \a4/a4/U5  ( .A(ts3[4]), .B(tc3[4]), .Y(n153) );
  OAI21X1 \a4/a4/U3  ( .A(n153), .B(n152), .C(n27), .Y(\a4/c5 ) );
  XOR2X1 \a4/a4/U2  ( .A(n152), .B(n153), .Y(s[4]) );
  XNOR2X1 \a4/a3/U5  ( .A(ts3[3]), .B(tc3[3]), .Y(n150) );
  OAI21X1 \a4/a3/U3  ( .A(n150), .B(n149), .C(n6), .Y(\a4/c4 ) );
  XOR2X1 \a4/a3/U2  ( .A(n149), .B(n150), .Y(s[3]) );
  XNOR2X1 \a4/a2/U5  ( .A(ts3[2]), .B(tc3[2]), .Y(n147) );
  OAI21X1 \a4/a2/U3  ( .A(n147), .B(n41), .C(n19), .Y(\a4/c3 ) );
  XOR2X1 \a4/a2/U2  ( .A(n41), .B(n147), .Y(s[2]) );
  XOR2X1 \a4/a1/U2  ( .A(n51), .B(n42), .Y(s[1]) );
  XOR2X1 \a4/a0/U2  ( .A(n146), .B(n2), .Y(s[0]) );
  XNOR2X1 \a3/s15/U5  ( .A(\a3/ts[5] ), .B(tc2[5]), .Y(n144) );
  OAI21X1 \a3/s15/U3  ( .A(n144), .B(n143), .C(n7), .Y(tc3[6]) );
  XOR2X1 \a3/s15/U2  ( .A(n143), .B(n144), .Y(ts3[5]) );
  XNOR2X1 \a3/s14/U5  ( .A(\a3/ts[4] ), .B(tc2[4]), .Y(n141) );
  OAI21X1 \a3/s14/U3  ( .A(n141), .B(n140), .C(n8), .Y(tc3[5]) );
  XOR2X1 \a3/s14/U2  ( .A(n140), .B(n141), .Y(ts3[4]) );
  XNOR2X1 \a3/s13/U5  ( .A(\a3/ts[3] ), .B(tc2[3]), .Y(n138) );
  OAI21X1 \a3/s13/U3  ( .A(n138), .B(n137), .C(n9), .Y(tc3[4]) );
  XOR2X1 \a3/s13/U2  ( .A(n137), .B(n138), .Y(ts3[3]) );
  XNOR2X1 \a3/s12/U5  ( .A(\a3/ts[2] ), .B(tc2[2]), .Y(n135) );
  OAI21X1 \a3/s12/U3  ( .A(n135), .B(n134), .C(n10), .Y(tc3[3]) );
  XOR2X1 \a3/s12/U2  ( .A(n134), .B(n135), .Y(ts3[2]) );
  XNOR2X1 \a3/s11/U5  ( .A(\a3/ts[1] ), .B(n56), .Y(n132) );
  OAI21X1 \a3/s11/U3  ( .A(n132), .B(n50), .C(n31), .Y(tc3[2]) );
  XNOR2X1 \a3/s05/U5  ( .A(ts1[5]), .B(tc1[5]), .Y(n130) );
  OAI21X1 \a3/s05/U3  ( .A(n130), .B(n49), .C(n11), .Y(\a3/tc[6] ) );
  XOR2X1 \a3/s05/U2  ( .A(n49), .B(n130), .Y(\a3/ts[5] ) );
  XNOR2X1 \a3/s04/U5  ( .A(ts1[4]), .B(tc1[4]), .Y(n128) );
  OAI21X1 \a3/s04/U3  ( .A(n128), .B(n48), .C(n12), .Y(\a3/tc[5] ) );
  XOR2X1 \a3/s04/U2  ( .A(n48), .B(n128), .Y(\a3/ts[4] ) );
  XNOR2X1 \a3/s03/U5  ( .A(ts1[3]), .B(tc1[3]), .Y(n126) );
  OAI21X1 \a3/s03/U3  ( .A(n126), .B(n47), .C(n13), .Y(\a3/tc[4] ) );
  XOR2X1 \a3/s03/U2  ( .A(n47), .B(n126), .Y(\a3/ts[3] ) );
  XNOR2X1 \a3/s02/U5  ( .A(ts1[2]), .B(tc1[2]), .Y(n124) );
  OAI21X1 \a3/s02/U3  ( .A(n124), .B(n44), .C(n14), .Y(\a3/tc[3] ) );
  XOR2X1 \a3/s02/U2  ( .A(n44), .B(n124), .Y(\a3/ts[2] ) );
  XNOR2X1 \a3/s01/U5  ( .A(ts1[1]), .B(n52), .Y(n122) );
  OAI21X1 \a3/s01/U3  ( .A(n122), .B(n43), .C(n15), .Y(\a3/tc[2] ) );
  XOR2X1 \a3/s01/U2  ( .A(n43), .B(n122), .Y(\a3/ts[1] ) );
  XNOR2X1 \a2/s16/U5  ( .A(\a2/ts[6] ), .B(h[6]), .Y(n121) );
  XOR2X1 \a2/s16/U2  ( .A(n120), .B(n121), .Y(\ts2[6] ) );
  XNOR2X1 \a2/s15/U5  ( .A(\a2/ts[5] ), .B(h[5]), .Y(n118) );
  OAI21X1 \a2/s15/U3  ( .A(n118), .B(n117), .C(n40), .Y(tc2[6]) );
  XNOR2X1 \a2/s14/U5  ( .A(\a2/ts[4] ), .B(h[4]), .Y(n115) );
  OAI21X1 \a2/s14/U3  ( .A(n115), .B(n114), .C(n18), .Y(tc2[5]) );
  XNOR2X1 \a2/s13/U5  ( .A(\a2/ts[3] ), .B(h[3]), .Y(n112) );
  OAI21X1 \a2/s13/U3  ( .A(n112), .B(n111), .C(n20), .Y(tc2[4]) );
  XNOR2X1 \a2/s12/U5  ( .A(\a2/ts[2] ), .B(h[2]), .Y(n109) );
  OAI21X1 \a2/s12/U3  ( .A(n109), .B(n108), .C(n22), .Y(tc2[3]) );
  XNOR2X1 \a2/s11/U5  ( .A(\a2/ts[1] ), .B(h[1]), .Y(n106) );
  OAI21X1 \a2/s11/U3  ( .A(n106), .B(n105), .C(n24), .Y(tc2[2]) );
  XNOR2X1 \a2/s05/U5  ( .A(e[5]), .B(f[5]), .Y(n103) );
  OAI21X1 \a2/s05/U3  ( .A(n103), .B(n102), .C(n29), .Y(\a2/tc[6] ) );
  XOR2X1 \a2/s05/U2  ( .A(n102), .B(n103), .Y(\a2/ts[5] ) );
  XNOR2X1 \a2/s04/U5  ( .A(e[4]), .B(f[4]), .Y(n100) );
  OAI21X1 \a2/s04/U3  ( .A(n100), .B(n99), .C(n26), .Y(\a2/tc[5] ) );
  XOR2X1 \a2/s04/U2  ( .A(n99), .B(n100), .Y(\a2/ts[4] ) );
  XNOR2X1 \a2/s03/U5  ( .A(e[3]), .B(f[3]), .Y(n97) );
  OAI21X1 \a2/s03/U3  ( .A(n97), .B(n96), .C(n32), .Y(\a2/tc[4] ) );
  XOR2X1 \a2/s03/U2  ( .A(n96), .B(n97), .Y(\a2/ts[3] ) );
  XNOR2X1 \a2/s02/U5  ( .A(e[2]), .B(f[2]), .Y(n94) );
  OAI21X1 \a2/s02/U3  ( .A(n94), .B(n93), .C(n34), .Y(\a2/tc[3] ) );
  XOR2X1 \a2/s02/U2  ( .A(n93), .B(n94), .Y(\a2/ts[2] ) );
  XNOR2X1 \a2/s01/U5  ( .A(e[1]), .B(f[1]), .Y(n91) );
  OAI21X1 \a2/s01/U3  ( .A(n91), .B(n90), .C(n36), .Y(\a2/tc[2] ) );
  XOR2X1 \a2/s01/U2  ( .A(n90), .B(n91), .Y(\a2/ts[1] ) );
  XNOR2X1 \a2/s00/U5  ( .A(e[0]), .B(f[0]), .Y(n88) );
  OAI21X1 \a2/s00/U3  ( .A(n88), .B(n87), .C(n38), .Y(\a2/tc[1] ) );
  XOR2X1 \a2/s00/U2  ( .A(n87), .B(n88), .Y(\a2/ts[0] ) );
  XNOR2X1 \a1/s15/U5  ( .A(\a1/ts[5] ), .B(d[5]), .Y(n85) );
  OAI21X1 \a1/s15/U3  ( .A(n85), .B(n84), .C(n17), .Y(tc1[6]) );
  XOR2X1 \a1/s15/U2  ( .A(n84), .B(n85), .Y(ts1[5]) );
  XNOR2X1 \a1/s14/U5  ( .A(\a1/ts[4] ), .B(d[4]), .Y(n82) );
  OAI21X1 \a1/s14/U3  ( .A(n82), .B(n81), .C(n16), .Y(tc1[5]) );
  XOR2X1 \a1/s14/U2  ( .A(n81), .B(n82), .Y(ts1[4]) );
  XNOR2X1 \a1/s13/U5  ( .A(\a1/ts[3] ), .B(d[3]), .Y(n79) );
  OAI21X1 \a1/s13/U3  ( .A(n79), .B(n78), .C(n21), .Y(tc1[4]) );
  XOR2X1 \a1/s13/U2  ( .A(n78), .B(n79), .Y(ts1[3]) );
  XNOR2X1 \a1/s12/U5  ( .A(\a1/ts[2] ), .B(d[2]), .Y(n76) );
  OAI21X1 \a1/s12/U3  ( .A(n76), .B(n75), .C(n23), .Y(tc1[3]) );
  XOR2X1 \a1/s12/U2  ( .A(n75), .B(n76), .Y(ts1[2]) );
  XNOR2X1 \a1/s11/U5  ( .A(\a1/ts[1] ), .B(d[1]), .Y(n73) );
  OAI21X1 \a1/s11/U3  ( .A(n73), .B(n72), .C(n25), .Y(tc1[2]) );
  XOR2X1 \a1/s11/U2  ( .A(n72), .B(n73), .Y(ts1[1]) );
  XNOR2X1 \a1/s05/U5  ( .A(a[5]), .B(b[5]), .Y(n70) );
  OAI21X1 \a1/s05/U3  ( .A(n70), .B(n69), .C(n30), .Y(\a1/tc[6] ) );
  XOR2X1 \a1/s05/U2  ( .A(n69), .B(n70), .Y(\a1/ts[5] ) );
  XNOR2X1 \a1/s04/U5  ( .A(a[4]), .B(b[4]), .Y(n67) );
  OAI21X1 \a1/s04/U3  ( .A(n67), .B(n66), .C(n28), .Y(\a1/tc[5] ) );
  XOR2X1 \a1/s04/U2  ( .A(n66), .B(n67), .Y(\a1/ts[4] ) );
  XNOR2X1 \a1/s03/U5  ( .A(a[3]), .B(b[3]), .Y(n64) );
  OAI21X1 \a1/s03/U3  ( .A(n64), .B(n63), .C(n33), .Y(\a1/tc[4] ) );
  XOR2X1 \a1/s03/U2  ( .A(n63), .B(n64), .Y(\a1/ts[3] ) );
  XNOR2X1 \a1/s02/U5  ( .A(a[2]), .B(b[2]), .Y(n61) );
  OAI21X1 \a1/s02/U3  ( .A(n61), .B(n60), .C(n35), .Y(\a1/tc[3] ) );
  XOR2X1 \a1/s02/U2  ( .A(n60), .B(n61), .Y(\a1/ts[2] ) );
  XNOR2X1 \a1/s01/U5  ( .A(a[1]), .B(b[1]), .Y(n58) );
  OAI21X1 \a1/s01/U3  ( .A(n58), .B(n57), .C(n37), .Y(\a1/tc[2] ) );
  XOR2X1 \a1/s01/U2  ( .A(n57), .B(n58), .Y(\a1/ts[1] ) );
  XNOR2X1 U1 ( .A(\a1/ts[0] ), .B(d[0]), .Y(n1) );
  XNOR2X1 U2 ( .A(n3), .B(n1), .Y(n2) );
  XNOR2X1 U3 ( .A(\a2/ts[0] ), .B(h[0]), .Y(n3) );
  AND2X1 U4 ( .A(ts3[5]), .B(tc3[5]), .Y(n157) );
  INVX1 U5 ( .A(n157), .Y(n4) );
  AND2X1 U6 ( .A(ts3[6]), .B(tc3[6]), .Y(n160) );
  INVX1 U7 ( .A(n160), .Y(n5) );
  AND2X1 U8 ( .A(ts3[3]), .B(tc3[3]), .Y(n151) );
  INVX1 U9 ( .A(n151), .Y(n6) );
  AND2X1 U10 ( .A(\a3/ts[5] ), .B(tc2[5]), .Y(n145) );
  INVX1 U11 ( .A(n145), .Y(n7) );
  AND2X1 U12 ( .A(\a3/ts[4] ), .B(tc2[4]), .Y(n142) );
  INVX1 U13 ( .A(n142), .Y(n8) );
  AND2X1 U14 ( .A(\a3/ts[3] ), .B(tc2[3]), .Y(n139) );
  INVX1 U15 ( .A(n139), .Y(n9) );
  AND2X1 U16 ( .A(\a3/ts[2] ), .B(tc2[2]), .Y(n136) );
  INVX1 U17 ( .A(n136), .Y(n10) );
  AND2X1 U18 ( .A(ts1[5]), .B(tc1[5]), .Y(n131) );
  INVX1 U19 ( .A(n131), .Y(n11) );
  AND2X1 U20 ( .A(ts1[4]), .B(tc1[4]), .Y(n129) );
  INVX1 U21 ( .A(n129), .Y(n12) );
  AND2X1 U22 ( .A(ts1[3]), .B(tc1[3]), .Y(n127) );
  INVX1 U23 ( .A(n127), .Y(n13) );
  AND2X1 U24 ( .A(ts1[2]), .B(tc1[2]), .Y(n125) );
  INVX1 U25 ( .A(n125), .Y(n14) );
  AND2X1 U26 ( .A(ts1[1]), .B(n52), .Y(n123) );
  INVX1 U27 ( .A(n123), .Y(n15) );
  AND2X1 U28 ( .A(\a1/ts[4] ), .B(d[4]), .Y(n83) );
  INVX1 U29 ( .A(n83), .Y(n16) );
  AND2X1 U30 ( .A(\a1/ts[5] ), .B(d[5]), .Y(n86) );
  INVX1 U31 ( .A(n86), .Y(n17) );
  AND2X1 U32 ( .A(\a2/ts[4] ), .B(h[4]), .Y(n116) );
  INVX1 U33 ( .A(n116), .Y(n18) );
  AND2X1 U34 ( .A(ts3[2]), .B(tc3[2]), .Y(n148) );
  INVX1 U35 ( .A(n148), .Y(n19) );
  AND2X1 U36 ( .A(\a2/ts[3] ), .B(h[3]), .Y(n113) );
  INVX1 U37 ( .A(n113), .Y(n20) );
  AND2X1 U38 ( .A(\a1/ts[3] ), .B(d[3]), .Y(n80) );
  INVX1 U39 ( .A(n80), .Y(n21) );
  AND2X1 U40 ( .A(\a2/ts[2] ), .B(h[2]), .Y(n110) );
  INVX1 U41 ( .A(n110), .Y(n22) );
  AND2X1 U42 ( .A(\a1/ts[2] ), .B(d[2]), .Y(n77) );
  INVX1 U43 ( .A(n77), .Y(n23) );
  AND2X1 U44 ( .A(\a2/ts[1] ), .B(h[1]), .Y(n107) );
  INVX1 U45 ( .A(n107), .Y(n24) );
  AND2X1 U46 ( .A(\a1/ts[1] ), .B(d[1]), .Y(n74) );
  INVX1 U47 ( .A(n74), .Y(n25) );
  AND2X1 U48 ( .A(e[4]), .B(f[4]), .Y(n101) );
  INVX1 U49 ( .A(n101), .Y(n26) );
  AND2X1 U50 ( .A(ts3[4]), .B(tc3[4]), .Y(n154) );
  INVX1 U51 ( .A(n154), .Y(n27) );
  AND2X1 U52 ( .A(a[4]), .B(b[4]), .Y(n68) );
  INVX1 U53 ( .A(n68), .Y(n28) );
  AND2X1 U54 ( .A(e[5]), .B(f[5]), .Y(n104) );
  INVX1 U55 ( .A(n104), .Y(n29) );
  AND2X1 U56 ( .A(a[5]), .B(b[5]), .Y(n71) );
  INVX1 U57 ( .A(n71), .Y(n30) );
  AND2X1 U58 ( .A(\a3/ts[1] ), .B(n56), .Y(n133) );
  INVX1 U59 ( .A(n133), .Y(n31) );
  AND2X1 U60 ( .A(e[3]), .B(f[3]), .Y(n98) );
  INVX1 U61 ( .A(n98), .Y(n32) );
  AND2X1 U62 ( .A(a[3]), .B(b[3]), .Y(n65) );
  INVX1 U63 ( .A(n65), .Y(n33) );
  AND2X1 U64 ( .A(e[2]), .B(f[2]), .Y(n95) );
  INVX1 U65 ( .A(n95), .Y(n34) );
  AND2X1 U66 ( .A(a[2]), .B(b[2]), .Y(n62) );
  INVX1 U67 ( .A(n62), .Y(n35) );
  AND2X1 U68 ( .A(e[1]), .B(f[1]), .Y(n92) );
  INVX1 U69 ( .A(n92), .Y(n36) );
  AND2X1 U70 ( .A(a[1]), .B(b[1]), .Y(n59) );
  INVX1 U71 ( .A(n59), .Y(n37) );
  AND2X1 U72 ( .A(e[0]), .B(f[0]), .Y(n89) );
  INVX1 U73 ( .A(n89), .Y(n38) );
  AND2X1 U74 ( .A(a[0]), .B(b[0]), .Y(\a1/s00/n3 ) );
  INVX1 U75 ( .A(\a1/s00/n3 ), .Y(n39) );
  AND2X1 U76 ( .A(\a2/ts[5] ), .B(h[5]), .Y(n119) );
  INVX1 U77 ( .A(n119), .Y(n40) );
  OR2X1 U78 ( .A(n42), .B(n51), .Y(n41) );
  XNOR2X1 U79 ( .A(n50), .B(n132), .Y(n42) );
  INVX1 U80 ( .A(\a4/c3 ), .Y(n149) );
  INVX1 U81 ( .A(\a4/c4 ), .Y(n152) );
  INVX1 U82 ( .A(\a4/c5 ), .Y(n155) );
  INVX1 U83 ( .A(\a4/c6 ), .Y(n158) );
  XNOR2X1 U84 ( .A(n105), .B(n106), .Y(n43) );
  XNOR2X1 U85 ( .A(n108), .B(n109), .Y(n44) );
  INVX1 U86 ( .A(\a3/tc[2] ), .Y(n134) );
  XOR2X1 U87 ( .A(\a3/tc[6] ), .B(n45), .Y(ts3[6]) );
  XOR2X1 U88 ( .A(\a3/ts[6] ), .B(tc2[6]), .Y(n45) );
  XOR2X1 U89 ( .A(\ts2[6] ), .B(n46), .Y(\a3/ts[6] ) );
  XOR2X1 U90 ( .A(ts1[6]), .B(tc1[6]), .Y(n46) );
  XNOR2X1 U91 ( .A(n111), .B(n112), .Y(n47) );
  XNOR2X1 U92 ( .A(n114), .B(n115), .Y(n48) );
  XNOR2X1 U93 ( .A(n117), .B(n118), .Y(n49) );
  INVX1 U94 ( .A(\a3/tc[3] ), .Y(n137) );
  INVX1 U95 ( .A(\a3/tc[4] ), .Y(n140) );
  INVX1 U96 ( .A(\a3/tc[5] ), .Y(n143) );
  OR2X1 U97 ( .A(n1), .B(n3), .Y(n50) );
  OR2X1 U98 ( .A(n2), .B(n146), .Y(n51) );
  INVX1 U99 ( .A(\a1/tc[1] ), .Y(n72) );
  INVX1 U100 ( .A(\a1/tc[2] ), .Y(n75) );
  AND2X1 U101 ( .A(\a1/ts[0] ), .B(d[0]), .Y(n52) );
  INVX1 U102 ( .A(c[0]), .Y(\a1/s00/n1 ) );
  INVX1 U103 ( .A(c[1]), .Y(n57) );
  INVX1 U104 ( .A(c[2]), .Y(n60) );
  XOR2X1 U105 ( .A(\a1/tc[6] ), .B(n53), .Y(ts1[6]) );
  XOR2X1 U106 ( .A(\a1/ts[6] ), .B(d[6]), .Y(n53) );
  XOR2X1 U107 ( .A(c[6]), .B(n54), .Y(\a1/ts[6] ) );
  XOR2X1 U108 ( .A(a[6]), .B(b[6]), .Y(n54) );
  XOR2X1 U109 ( .A(g[6]), .B(n55), .Y(\a2/ts[6] ) );
  XOR2X1 U110 ( .A(e[6]), .B(f[6]), .Y(n55) );
  INVX1 U111 ( .A(\a2/tc[1] ), .Y(n105) );
  INVX1 U112 ( .A(\a2/tc[2] ), .Y(n108) );
  INVX1 U113 ( .A(\a1/tc[3] ), .Y(n78) );
  INVX1 U114 ( .A(\a2/tc[3] ), .Y(n111) );
  INVX1 U115 ( .A(\a1/tc[4] ), .Y(n81) );
  INVX1 U116 ( .A(\a2/tc[4] ), .Y(n114) );
  INVX1 U117 ( .A(\a2/tc[5] ), .Y(n117) );
  INVX1 U118 ( .A(\a1/tc[5] ), .Y(n84) );
  INVX1 U119 ( .A(\a2/tc[6] ), .Y(n120) );
  AND2X1 U120 ( .A(\a2/ts[0] ), .B(h[0]), .Y(n56) );
  INVX1 U121 ( .A(g[0]), .Y(n87) );
  INVX1 U122 ( .A(g[1]), .Y(n90) );
  INVX1 U123 ( .A(g[2]), .Y(n93) );
  INVX1 U124 ( .A(c[3]), .Y(n63) );
  INVX1 U125 ( .A(g[3]), .Y(n96) );
  INVX1 U126 ( .A(c[4]), .Y(n66) );
  INVX1 U127 ( .A(g[4]), .Y(n99) );
  INVX1 U128 ( .A(g[5]), .Y(n102) );
  INVX1 U129 ( .A(c[5]), .Y(n69) );
  INVX1 U130 ( .A(ci), .Y(n146) );
endmodule

